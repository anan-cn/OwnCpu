----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:48:06 03/13/2013 
-- Design Name: 
-- Module Name:    InstrMem32bit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstrMem32bit is
    Port ( address : in  STD_LOGIC_VECTOR (31 downto 0);
           Instr : out  STD_LOGIC_VECTOR (31 downto 0));
end InstrMem32bit;


architecture Behavioral of InstrMem32bit is

type ARRAY_256 is ARRAY (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
signal MemContent: ARRAY_256 :=	(	X"00000063",X"0000007c",X"00000077",X"0000007b",X"000000f2",X"0000006b",X"0000006f",X"000000c5",X"00000002",X"00000001",X"00000067",X"0000002b",X"000000fe",X"000000d7",X"000000ab",X"00000076",
											X"000000ca",X"00000082",X"000000c9",X"0000007d",X"000000fa",X"00000059",X"00000047",X"000000f0",X"000000ad",X"000000d4",X"000000a2",X"000000af",X"0000009c",X"000000a4",X"00000072",X"000000c0",
											X"000000b7",X"000000fd",X"00000093",X"00000026",X"00000036",X"0000003f",X"000000f7",X"000000cc",X"00000034",X"000000a5",X"000000e5",X"000000f1",X"00000071",X"000000d8",X"00000031",X"00000015",
											X"00000004",X"000000c7",X"00000023",X"000000c3",X"00000018",X"00000096",X"00000005",X"0000009a",X"00000007",X"00000012",X"00000080",X"000000e2",X"000000eb",X"00000027",X"000000b2",X"00000075",
											X"00000009",X"00000083",X"0000002c",X"0000001a",X"0000001b",X"0000006e",X"0000005a",X"000000a0",X"00000052",X"0000003b",X"000000d6",X"000000b3",X"00000029",X"000000e3",X"0000002f",X"00000084",
											X"00000053",X"000000d1",X"00000000",X"000000ed",X"00000020",X"000000fc",X"000000b1",X"0000005b",X"0000006a",X"000000cb",X"000000be",X"00000039",X"0000004a",X"0000004c",X"00000058",X"000000cf",
											X"000000d0",X"000000ef",X"000000aa",X"000000fb",X"00000043",X"0000004d",X"00000033",X"00000085",X"00000045",X"000000f9",X"00000002",X"0000007f",X"00000050",X"0000003c",X"0000009f",X"000000a8",
											X"00000051",X"000000a3",X"00000040",X"0000008f",X"00000092",X"0000009d",X"00000038",X"000000f5",X"000000bc",X"000000b6",X"000000da",X"00000021",X"00000010",X"000000ff",X"000000f3",X"000000d2",
											X"000000cd",X"0000000c",X"00000013",X"000000ec",X"0000005f",X"00000097",X"00000044",X"00000017",X"000000c4",X"000000a7",X"0000007e",X"0000003d",X"00000064",X"0000005d",X"00000019",X"00000073",
											X"00000060",X"00000081",X"0000004f",X"000000dc",X"00000022",X"0000002a",X"00000090",X"00000088",X"00000046",X"000000ee",X"000000b8",X"00000014",X"000000de",X"0000005e",X"0000000b",X"000000db",
											X"000000e0",X"00000032",X"0000003a",X"0000000a",X"00000049",X"00000006",X"00000024",X"0000005c",X"000000c2",X"000000d3",X"000000ac",X"00000062",X"00000091",X"00000095",X"000000e4",X"00000079",
											X"000000e7",X"000000c8",X"00000037",X"0000006d",X"0000008d",X"000000d5",X"0000004e",X"000000a9",X"0000006c",X"00000056",X"000000f4",X"000000ea",X"00000065",X"0000007a",X"000000ae",X"00000008",
											X"000000ba",X"00000078",X"00000025",X"0000002e",X"0000001c",X"000000a6",X"000000b4",X"000000c6",X"000000e8",X"000000dd",X"00000074",X"0000001f",X"0000004b",X"000000bd",X"0000008b",X"0000008a",
											X"00000070",X"0000003e",X"000000b5",X"00000066",X"00000048",X"00000003",X"000000f6",X"0000000e",X"00000061",X"00000035",X"00000057",X"000000b9",X"00000086",X"000000c1",X"0000001d",X"0000009e",
											X"000000e1",X"000000f8",X"00000098",X"00000011",X"00000069",X"000000d9",X"0000008e",X"00000094",X"0000009b",X"0000001e",X"00000087",X"000000e9",X"000000ce",X"00000055",X"00000028",X"000000df",
											X"0000008c",X"000000a1",X"00000089",X"0000000d",X"000000bf",X"000000e6",X"00000042",X"00000068",X"00000041",X"00000099",X"0000002d",X"0000000f",X"000000b0",X"00000054",X"000000bb",X"00000016"	);

begin

--Instr<=MemContent(to_integer(unsigned(address) srl 2) );
Instr <= MemContent(to_integer(unsigned(address(31 downto 2))));

end Behavioral;

